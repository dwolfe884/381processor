library IEEE;
use IEEE.std_logic_1164.all;

entity tb_mux31t1 is
  generic(N : integer := 32;
          gCLK_HPER   : time := 50 ns);
end tb_mux31t1;

architecture behavior of tb_mux31t1 is
  
  -- Calculate the clock period as twice the half-period
  constant cCLK_PER  : time := gCLK_HPER * 2;


  component mux31t1
    port(i_0          : in std_logic_vector(31 downto 0);
       i_1          : in std_logic_vector(31 downto 0); 
       i_2          : in std_logic_vector(31 downto 0);
       i_3          : in std_logic_vector(31 downto 0);
       i_4          : in std_logic_vector(31 downto 0);
       i_5          : in std_logic_vector(31 downto 0);
       i_6          : in std_logic_vector(31 downto 0);
       i_7          : in std_logic_vector(31 downto 0);
       i_8          : in std_logic_vector(31 downto 0);
       i_9          : in std_logic_vector(31 downto 0);
       i_10          : in std_logic_vector(31 downto 0);
       i_11          : in std_logic_vector(31 downto 0);
       i_12          : in std_logic_vector(31 downto 0);
       i_13          : in std_logic_vector(31 downto 0);
       i_14          : in std_logic_vector(31 downto 0);
       i_15          : in std_logic_vector(31 downto 0);
       i_16          : in std_logic_vector(31 downto 0);
       i_17          : in std_logic_vector(31 downto 0);
       i_18          : in std_logic_vector(31 downto 0);
       i_19          : in std_logic_vector(31 downto 0);
       i_20          : in std_logic_vector(31 downto 0);
       i_21          : in std_logic_vector(31 downto 0);
       i_22          : in std_logic_vector(31 downto 0);
       i_23          : in std_logic_vector(31 downto 0);
       i_24          : in std_logic_vector(31 downto 0);
       i_25          : in std_logic_vector(31 downto 0);
       i_26          : in std_logic_vector(31 downto 0);
       i_27          : in std_logic_vector(31 downto 0);
       i_28          : in std_logic_vector(31 downto 0);
       i_29          : in std_logic_vector(31 downto 0);
       i_30          : in std_logic_vector(31 downto 0);
       i_31          : in std_logic_vector(31 downto 0);
       i_s	     : in std_logic_vector(4 downto 0);
       o_out          : out std_logic_vector(31 downto 0));

  end component;

  -- Temporary signals to connect to the dff component.
  signal s_0,s_1,s_2,s_3,s_4,s_5,s_6,s_7,s_8,s_9,s_10,s_11,s_12,s_13,s_14,s_15,s_16,s_17,s_18,s_19,s_20,s_21,s_22,s_23,s_24,s_25,s_26,s_27,s_28,s_29,s_30,s_31 : std_logic_vector(31 downto 0) := x"00000000";
  signal s_s : std_logic_vector(4 downto 0):= "00000"; 
  signal s_out : std_logic_vector(31 downto 0);

begin

  DUT: mux31t1 
  port map(i_0   => s_0,
	i_1   => s_1,
	i_2   => s_2,
	i_3   => s_3,
	i_4   => s_4,
	i_5   => s_5,
	i_6   => s_6,
	i_7   => s_7,
	i_8   => s_8,
	i_9   => s_9,
	i_10   => s_10,
	i_11   => s_11,
	i_12   => s_12,
	i_13   => s_13,
	i_14   => s_14,
	i_15   => s_15,
	i_16   => s_16,
	i_17   => s_17,
	i_18   => s_18,
	i_19   => s_19,
	i_20   => s_20,
	i_21   => s_21,
	i_22   => s_22,
	i_23   => s_23,
	i_24   => s_24,
	i_25   => s_25,
	i_26   => s_26,
	i_27   => s_27,
	i_28   => s_28,
	i_29   => s_29,
	i_30   => s_30,
	i_31   => s_31,
	   i_s    => s_s,
           o_out   => s_out);

  -- Testbench process  
  P_TB: process
  begin
    s_0   <= x"00000000";
    s_1   <= x"00000001";
    s_2   <= x"00000002";
    s_3   <= x"00000003";
    s_4   <= x"00000004";
    s_5   <= x"00000005";
    s_6   <= x"00000006";
    s_7   <= x"00000007";

    -- Reset the FF
    s_s   <= "00000";
    wait for cCLK_PER;
    s_s   <= "00001";
    wait for cCLK_PER;
    s_s   <= "00010";
    wait for cCLK_PER;
    s_s   <= "00011";
    wait for cCLK_PER;
    s_s   <= "00100";
    wait for cCLK_PER;
    s_s   <= "00101";
    wait for cCLK_PER;
    s_s   <= "00110";
    wait for cCLK_PER;
    s_s   <= "00111";
    wait for cCLK_PER;
    s_s   <= "01000";
    wait for cCLK_PER;
    s_s   <= "01001";
    wait for cCLK_PER;
    s_s   <= "01011";
    wait for cCLK_PER;
    s_s   <= "01100";
    wait for cCLK_PER;
    s_s   <= "01101";
    wait for cCLK_PER;
    s_s   <= "01110";
    wait for cCLK_PER;
    s_s   <= "01111";
    wait for cCLK_PER;
  end process;
  
end behavior;