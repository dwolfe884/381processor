library IEEE;
use IEEE.std_logic_1164.all;

entity cu is

  port(i_op     : in std_logic_vector(5 downto 0);
       i_func   : in std_logic_vector(5 downto 0);
       aluControl   : out std_logic_vector(3 downto 0);
       b        : out std_logic;
       j	: out std_logic;
       jr	: out std_logic;
       jal	: out std_logic;
       memRead  : out std_logic;
       memToReg : out std_logic;
       memWrite : out std_logic;
       aluSrc   : out std_logic;
       regWrite : out std_logic;
       sign_ext	: out std_logic;
       regDst   : out std_logic;
       vsig	: out std_logic;
       halt	: out std_logic);
       
end cu;

architecture mixed of cu is
begin
process(i_op, i_func)
begin
    jr <= '0';
    jal <= '0';
    vsig <= '1';
    halt <= '0';
    if (i_op = "001000") then --addi
	aluControl <= "0000";
	regDst <= '0';
        aluSrc <= '1';
        memToReg <= '0';
        regWrite <= '1';
        memRead <= '0';
        memWrite <= '0';
	sign_ext <= '1';
        b <= '0';
	j <= '0';
    elsif i_op = "010100" then --halt
	aluControl <= "0000";
	regDst <= '0';
        aluSrc <= '0';
        memToReg <= '0';
        regWrite <= '0';
        memRead <= '0';
        memWrite <= '0';
	sign_ext <= '0';
        b <= '0';
	j <= '0';
	halt <= '1';
    elsif i_op = "001001" then --addiu
	aluControl <= "0000";
	regDst <= '0';
        aluSrc <= '1';
        memToReg <= '0';
        regWrite <= '1';
        memRead <= '0';
        memWrite <= '0';
	sign_ext <= '1';
        b <= '0';
	j <= '0';
	vsig <= '0';
    elsif i_op = "000000" then 
        if i_func = "100000" then --add
            aluControl <= "0000";
            regDst <= '1';
            aluSrc <= '0';
            memToReg <= '0';
            regWrite <= '1';
            memRead <= '0';
            memWrite <= '0';
	    sign_ext <= '1';
            b <= '0';
            j <= '0';
	elsif i_func = "100001" then --addu
            aluControl <= "0000";
            regDst <= '1';
            aluSrc <= '0';
            memToReg <= '0';
            regWrite <= '1';
            memRead <= '0';
            memWrite <= '0';
	    sign_ext <= '0';
            b <= '0';
	    j <= '0';
	    vsig <= '0';
	elsif i_func = "100010" then --sub
            aluControl <= "1000";
            regDst <= '1';
            aluSrc <= '0';
            memToReg <= '0';
            regWrite <= '1';
            memRead <= '0';
            memWrite <= '0';
	    sign_ext <= '1';
            b <= '0';
	    j <= '0';
	elsif i_func = "100011" then --subu
            aluControl <= "1000";
            regDst <= '1';
            aluSrc <= '0';
            memToReg <= '0';
            regWrite <= '1';
            memRead <= '0';
            memWrite <= '0';
	    sign_ext <= '0';
            b <= '0';
	    j <= '0';
	    vsig <= '0';
	elsif i_func = "100100" then --and
            aluControl <= "0001";
            regDst <= '1';
            aluSrc <= '0';
            memToReg <= '0';
            regWrite <= '1';
            memRead <= '0';
            memWrite <= '0';
	    sign_ext <= '0';
            b <= '0';
	    j <= '0';
	elsif i_func = "100101" then --or
            aluControl <= "1011";
            regDst <= '1';
            aluSrc <= '0';
            memToReg <= '0';
            regWrite <= '1';
            memRead <= '0';
            memWrite <= '0';
	    sign_ext <= '0';
            b <= '0';
	    j <= '0';
	elsif i_func = "100110" then --xor
            aluControl <= "1001";
            regDst <= '1';
            aluSrc <= '0';
            memToReg <= '0';
            regWrite <= '1';
            memRead <= '0';
            memWrite <= '0';
	    sign_ext <= '0';
            b <= '0';
	    j <= '0';
	elsif i_func = "100111" then --nor
            aluControl <= "1100";
            regDst <= '1';
            aluSrc <= '0';
            memToReg <= '0';
            regWrite <= '1';
            memRead <= '0';
            memWrite <= '0';
	    sign_ext <= '0';
            b <= '0';
	    j <= '0';
	elsif i_func = "000000" then --sll
            aluControl <= "1110";
            regDst <= '1';
            aluSrc <= '0';
            memToReg <= '0';
            regWrite <= '1';
            memRead <= '0';
            memWrite <= '0';
	    sign_ext <= '0';
            b <= '0';
	    j <= '0';
	elsif i_func = "000010" then --srl
            aluControl <= "1111";
            regDst <= '1';
            aluSrc <= '0';
            memToReg <= '0';
            regWrite <= '1';
            memRead <= '0';
            memWrite <= '0';
	    sign_ext <= '0';
            b <= '0';
	    j <= '0';
	elsif i_func = "000011" then --sra
            aluControl <= "0110";
            regDst <= '1';
            aluSrc <= '0';
            memToReg <= '0';
            regWrite <= '1';
            memRead <= '0';
            memWrite <= '0';
	    sign_ext <= '0';
            b <= '0';
	    j <= '0';
	elsif i_func = "101010" then --slt
            aluControl <= "1010";
            regDst <= '1';
            aluSrc <= '0';
            memToReg <= '0';
            regWrite <= '1';
            memRead <= '0';
            memWrite <= '0';
	    sign_ext <= '0';
            b <= '0';
	    j <= '0';
	    vsig <= '0';
	elsif i_func = "001000" then --jr
            aluControl <= "0000";
            regDst <= '0';
            aluSrc <= '0';
            memToReg <= '0';
            regWrite <= '0';
            memRead <= '0';
            memWrite <= '0';
	    sign_ext <= '0';
	    jr <= '1';
            b <= '0';
	    j <= '0';
	else
	    aluControl <= "0000";
            regDst <= '0';
            aluSrc <= '0';
            memToReg <= '0';
            regWrite <= '0';
            memRead <= '0';
            memWrite <= '0';
	    sign_ext <= '0';
	    jr <= '0';
            b <= '0';
	    j <= '0';
        end if;
    elsif i_op = "100011" then --lw
	aluControl <= "0000";
	regDst <= '0';
        aluSrc <= '1';
        memToReg <= '1';
        regWrite <= '1';
        memRead <= '0';
        memWrite <= '0';
	sign_ext <= '1';
        b <= '0';
	j <= '0';
    elsif i_op = "101011" then --sw
	aluControl <= "0000";
	regDst <= '0';
        aluSrc <= '1';
        memToReg <= '0';
        regWrite <= '0';
        memRead <= '0';
        memWrite <= '1';
	sign_ext <= '1';
        b <= '0';
	j <= '0';
    elsif i_op = "001111" then --lui
	aluControl <= "0011";
	regDst <= '0';
        aluSrc <= '1';
        memToReg <= '0';
        regWrite <= '1';
        memRead <= '0';
        memWrite <= '0';
	sign_ext <= '1';
        b <= '0';
	j <= '0';
    elsif i_op = "001100" then --andi
            aluControl <= "0001";
            regDst <= '0';
            aluSrc <= '1';
            memToReg <= '0';
            regWrite <= '1';
            memRead <= '0';
            memWrite <= '0';
	    sign_ext <= '0';
            b <= '0';
	    j <= '0';
    elsif i_op = "001101" then --ori
	aluControl <= "1011";
            regDst <= '0';
            aluSrc <= '1';
            memToReg <= '0';
            regWrite <= '1';
            memRead <= '0';
            memWrite <= '0';
	    sign_ext <= '0';
            b <= '0';
	    j <= '0';
    elsif i_op = "001110" then --xori
	aluControl <= "1001";
            regDst <= '0';
            aluSrc <= '1';
            memToReg <= '0';
            regWrite <= '1';
            memRead <= '0';
            memWrite <= '0';
	    sign_ext <= '0';
            b <= '0';
	    j <= '0';
    elsif i_op = "001010" then --slti
	aluControl <= "1010";
            regDst <= '0';
            aluSrc <= '1';
            memToReg <= '0';
            regWrite <= '1';
            memRead <= '0';
            memWrite <= '0';
	    sign_ext <= '1';
            b <= '0';
	    j <= '0';
    elsif i_op = "000100" then --beq
	aluControl <= "1000";
            regDst <= '0';
            aluSrc <= '0';
            memToReg <= '0';
            regWrite <= '0';
            memRead <= '0';
            memWrite <= '0';
	    sign_ext <= '0';
            b <= '1';
	    j <= '0';
    elsif i_op = "000101" then --bne
	aluControl <= "0101";
            regDst <= '0';
            aluSrc <= '0';
            memToReg <= '0';
            regWrite <= '0';
            memRead <= '0';
            memWrite <= '0';
	    sign_ext <= '1';
            b <= '1';
	    j <= '0';
    elsif i_op = "000010" then --j
	aluControl <= "0000";
            regDst <= '0';
            aluSrc <= '0';
            memToReg <= '0';
            regWrite <= '0';
            memRead <= '0';
            memWrite <= '0';
	    sign_ext <= '0';
            b <= '0';
	    j <= '1';
	    jal <= '0';
    elsif i_op = "000011" then --jal
	aluControl <= "0000";
            regDst <= '0';
            aluSrc <= '0';
            memToReg <= '0';
            regWrite <= '1';
            memRead <= '0';
            memWrite <= '0';
	    sign_ext <= '0';
            b <= '0';
	    j <= '1';
	    jal <= '1';
    elsif i_op = "011111" then --repl.qb
	aluControl <= "0100";
            regDst <= '1';
            aluSrc <= '0';
            memToReg <= '0';
            regWrite <= '1';
            memRead <= '0';
            memWrite <= '0';
	    sign_ext <= '0';
            b <= '0';
	    j <= '0';
	    jal <= '0';
    else
	    aluControl <= "0000";
            regDst <= '0';
            aluSrc <= '0';
            memToReg <= '0';
            regWrite <= '0';
            memRead <= '0';
            memWrite <= '0';
	    sign_ext <= '0';
	    jr <= '0';
            b <= '0';
	    j <= '0';
    end if;
    end process;
  
end mixed;
